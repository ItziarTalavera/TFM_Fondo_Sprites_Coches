----------------------------------------------------------------------------------
--                            Tabla de nombre                                   --
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
library WORK;
use WORK.VGA_PKG.ALL;

entity tabla_nombre is
	port (
	--Puertos de entrada
	clk          	  : in std_logic;
	dir_tabla_nombre  : in std_logic_vector(10-1 downto 0); --960 posiciones de memoria
 	--Puertos de salida
	dato_tabla_nombre : out std_logic_vector(8-1 downto 0)
);
end tabla_nombre;

architecture behavioral of tabla_nombre is

signal dir_int_img : natural range 0 to 2**10-1;
type img is array (natural range<>) of std_logic_vector(8-1 downto 0);
constant title : img := (
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000000",
	"00000000",
	"00000000",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000000",
	"00000000",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000000",
	"00000000",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000000",
	"00000000",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000000",
	"00000000",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000000",
	"00000000",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000000",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000000",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000000",
	"00000000",
	"00000000",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000000",
	"00000000",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000000",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000000",
	"00000000",
	"00000000",
	"00000010",
	"00000000",
	"00000000",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000000",
	"00000000",
	"00000010",
	"00000010",
	"00000010",
	"00000000",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000000",
	"00000000",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000000",
	"00000000",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000000",
	"00000010",
	"00000010",
	"00000010",
	"00000000",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000000",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000000",
	"00000000",
	"00000010",
	"00000010",
	"00000000",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000000",
	"00000000",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000000",
	"00000000",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000000",
	"00000010",
	"00000010",
	"00000000",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000000",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000000",
	"00000010",
	"00000010",
	"00000000",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000000",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000000",
	"00000000",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000000",
	"00000010",
	"00000010",
	"00000000",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000000",
	"00000000",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000000",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000000",
	"00000000",
	"00000010",
	"00000010",
	"00000000",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000000",
	"00000000",
	"00000000",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000000",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000000",
	"00000000",
	"00000000",
	"00000010",
	"00000010",
	"00000010",
	"00000000",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000000",
	"00000000",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000000",
	"00000011",
	"00000011",
	"00000011",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000000",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000000",
	"00000000",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000000",
	"00000011",
	"00000011",
	"00000011",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000000",
	"00000000",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000000",
	"00000000",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000000",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000000",
	"00000000",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000000",
	"00000000",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000000",
	"00000000",
	"00000010",
	"00000010",
	"00000010",
	"00000000",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000000",
	"00000000",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000000",
	"00000000",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000000",
	"00000010",
	"00000010",
	"00000010",
	"00000000",
	"00000000",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000000",
	"00000000",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000000",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000000",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000000",
	"00000000",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000000",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000000",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000000",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000000",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000000",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000000",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000001",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000000",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000000",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000001",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000000",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000000",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000001",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000000",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000000",
	"00000000",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000001",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000000",
	"00000000",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000000",
	"00000000",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000001",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000011",
	"00000000",
	"00000000",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010",
	"00000010"
);

begin

dir_int_img <= to_integer(unsigned(dir_tabla_nombre));

P_img: process (clk)
begin
	if clk'event and clk='1' then
		dato_tabla_nombre <= title(dir_int_img);
	end if;
end process;

end behavioral;